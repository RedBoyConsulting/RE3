��%�5�E�T�d�t���������������������������������������������������������������������������������� �  `     ��   @  ����x��@�  ��������n��@�  �������� n@T <<      �����   � � � �  _@O9==      �����   � � � �  _@P9>>      �����   � � � �  x@Q9??      �����   � � � �  x@S9@@      �����  
 � � � �  i@Q9AA      �����   � � � �  n@`9BB      �����   � � � �  x@[ CC      �����   � � � �  x@\ DD      �����   � � � �  x@^ EE      �����  	 � � � �  x@i;FF      �����   � � � �  d@iGG      �����   � � � �  U@kHH      �����   � � � �  d@kII      �����   � � � �  x@jJJ      �����   � � � �  x@gKK      �����   � � � �   Z@Z9<<      �����  � � � �    ~�n2
�~&�"�N �"
` $a 4�D�@I  �   �      ��   @  ����x��@�  ��������   @S;;;      �����   � � � �   x@Z9<<      �����   � � � �   x@[9==      �����   � � � �   P@J >>      �����   � � � �   x@]9??      �����   � � � �    ���(	    
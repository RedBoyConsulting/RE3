��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��� �  �     ��   @  ����x��@�  ��������x��@�  �������� P@V'<<      �����  	 � � � �  K@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  s@a'GG      �����   � � � �  n@b'HH      �����   � � � �  n@c'II      �����   � � � �  }@d'JJ      �����   � � � �  i@U <<      �����  � � � �  s@U ==      �����  � � � �  s@V >>      �����  � � � �  x@W ??      �����  � � � �    8�	.,b�V�|r#�&$-2�8:p=    
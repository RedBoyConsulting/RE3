 � %� 5� E� S�? c�? s�? ��? ��? ��?���� � ������ �g  �� �    �     ��   @  ����d��@�  ��������  i@M9;;      �����   � � � �   x@N9<<      �����  	 � � � �   x@O9==      �����  
 � � � �   n@P9>>      �����   � � � �   n@W ??      �����   � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �   d@^'DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   A@T HH      �����M   � � � �    Z �<���J
��    
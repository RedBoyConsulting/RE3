��%�4�D�T�d�t�������������������$�����������������������������������������������������0Z �  �     ��   @  ������@�  ��������x��@�  ��������  d@T <<      �����   � � � �   @Vm==      �����   � � � �   x@V >>      �����   � � � �   n@]9??      �����   � � � �   n@c;@@      �����   � � � �   d@Y AA      �����   � � � �   }@XmBB      �����   � � � �   x@a9CC      �����   � � � �   @^'DD      �����   � � � �   x@a>EE      �����   � � � �   n@d9FF      �����  	 � � � �   n@e9GG      �����   � � � �   A@] HH      �����   � � � �   s@c'II      �����  
 � � � �   n@m'JJ      �����   � � � �   A@]9KK      �����   � � � �   Z@\9<<      �����  � � � �   Z@U ==      �����  � � � �   n@W >>      �����  � � � �    �@��F
�*��Hpf�!$#|%F+        
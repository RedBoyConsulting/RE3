�������������� S�? c�? s�? ��?���� ��?�������� ������ �������&   �     ��  	 @  ����d��@�  ��������  d B9<<      �����   � � � �   dB9<<      �����   � � � �   d B9<<      �����   � � � �   dB9<<      �����   � � � �    @S;??      �����   � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �    @S;DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   @Z9HH      �����  	 � � � �    Z �<��-�U�d            
��+�5�A�T�k�|������������������������������������������������������������������������������������L 0       ��   @  ����d��@�  �������� Z@N9<<      �����   � � � �  d@M9==      �����   � � � �  @Cm>>      �����_   � � � �  @DF??      �����_   � � � �  s@U9@@      �����   � � � �  x@DFAA      �����_   � � � �  @MXBB      �����_   � � � �  @NZCC      �����_   � � � �  d@_9DD      �����   � � � �  <@X9EE      �����  
 � � � �  P@b FF      �����   � � � �  d@_ GG      �����   � � � �  A@T HH      �����   � � � �  F@U II      �����   � � � �  P@X JJ      �����   � � � �   $@`����&� ~!�"$�%�)  
���������������� S�? c�? s�? ��?�������� �� ��@� ����������0@ P  0     ��   @  ����d��@�  ��������  Z@H <<      �����   � � � �   Z@H <<      �����   � � � �    @S;>>      �����   � � � �    @S;??      �����   � � � �    @S;??      �����   � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �    @S;DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   2@T HH      �����   � � � �   Z@U II      �����   � � � �   n@\9JJ      �����   � � � �    Z �<�&nv�"$(    
��%�5�E�T�d�u�������������������$���S�3�A�d�t���������������P� �  @     ��    @  ����x��@�  ��������s��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  x@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �  P@V'<<      �����  � � � �  K@W'==      ����� 	 � � � �  @Tm>>      ����� 
 � � � �  _@U9??      �����  � � � �  _@X @@      �����  � � � �  _@S9AA      �����  � � � �    @S;BB      �����  � � � �    @S;CC      �����  � � � �  n@[ DD      �����  � � � �  @\ EE      �����  � � � �  @[mFF      �����  � � � �  n@c GG      �����  � � � �  _@g9HH      �����  � � � �  i@g9II      �����  � � � �  i@h9JJ      �����  � � � �  i@i9KK      �����  � � � �    8�TV
N�`�4���t�L#T'*~.�/p27T8:�;�>�?  
B` 5` A�Ua ea ua ���������������������������������������������������������������������������������������������������������x  @  0     ��   @  ����d��@�  ��������   @S;;;      �����   � � � �   _@H <<      �����   � � � �  _@H <<      �����   � � � �  _@I ==      �����   � � � �  F@J >>      �����   � � � �  Z@Q9??      �����   � � � �  @R9@@      �����   � � � �  Z@M AA      �����   � � � �    ��<d�
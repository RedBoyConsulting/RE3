B` U` ����e` ua ������������������������������������������������B5���������������������������������������������������������py  @  0     ��   @  ����d��@�  ��������   @S;;;      �����   � � � �   x@H <<      �����   � � � �  x@H <<      �����   � � � �   n@M>==      �����   � � � �  n@M>==      �����   � � � �  n@J >>      �����   � � � �  x@K ??      �����   � � � �  x@L @@      �����   � � � �    N2��.  
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�� �  P     ��   @  ����i��@�  ��������i��@�  ��������  �� �  ��������  A@Z9<<      �����   � � � �  7@[9==      �����   � � � �  @Tm>>      �����   � � � �  s@Q9??      �����  	 � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@a9CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@f9GG      �����  
 � � � �  i@f9HH      �����   � � � �  _@h9II      �����   � � � �  n@h9JJ      �����   � � � �  _@Z9<<      �����  � � � �  i@[9==      �����  � � � �  i@\9>>      �����  � � � �  U@]9??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    822���
�F���vr *$|%F)�-<2b3    
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@a'GG      �����   � � � �  d@c'HH      �����   � � � �  d@b'II      �����   � � � �  d@d'JJ      �����   � � � �  Z@Z9<<      �����  � � � �  d@[9==      �����  � � � �  _@\9>>      �����  � � � �  U@]9??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b�~�*�$�%$)v*@.�267    
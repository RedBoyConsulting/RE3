��%�5�E�T�d�u�������������������$���������������������������������������������`� P        ��   @  ����x��@�  ��������d��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  x@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����  
 � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����  	 � � � �  x@N9<<      �����  � � � �  P@O9==      �����  � � � �  A@V >>      �����  � � � �  _@g9HH      �����  � � � �  d@j9II      �����  � � � �  Z@i9JJ      �����  � � � �  i@i9KK      �����  � � � �    8�TV
�D�6��z�!�"b$�'.,>/�2,6
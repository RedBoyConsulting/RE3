��$���S�3�A�d�t��������������������������������������������������������������������������������* p  @     ��   @  ����i��@�  ��������  �� �  ��������  A@Z9<<      �����   � � � �  7@[9==      �����   � � � �  @Tm>>      �����   � � � �  s@Q9??      �����  	 � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@a9CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@f9GG      �����  
 � � � �  i@f9HH      �����   � � � �  _@h9II      �����   � � � �  n@h9JJ      �����   � � � �    822���
�F���vr *$P%            
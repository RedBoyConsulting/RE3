 � %� 5� E� S�? c�? s�? ��? ��? ��? ��? � ��@�� �g ����P�  0       ��   @  ����d��@�  ��������  }@M9;;      �����   � � � �   n@N9<<      �����  	 � � � �   i@O9==      �����  
 � � � �   i@Tm>>      �����   � � � �   }C]9??      �����   � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �   d@^'DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   n@d>HH      �����   � � � �  n@d>HH      �����   � � � �    Z �<��(����    
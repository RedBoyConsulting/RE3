��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��x �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@e9GG      �����   � � � �  d@f9HH      �����   � � � �  d@g9II      �����   � � � �  d@h9JJ      �����   � � � �  Z@Z9<<      �����  � � � �  d@[9==      �����  � � � �  _@\9>>      �����  � � � �  U@]9??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b��X"d$\%h',/    
��%�5�E�T�d�t����������������������������������������������������������������������������������G `  0     ��   @  ����x��@�  �������� n@T <<      �����   � � � �  _@O9==      �����   � � � �  _@P9>>      �����   � � � �  x@Q9??      �����   � � � �  x@S9@@      �����   � � � �  i@Q9AA      �����   � � � �  n@`9BB      �����   � � � �  x@[ CC      �����   � � � �  x@\ DD      �����   � � � �  x@^ EE      �����   � � � �  x@i;FF      �����   � � � �  d@e9GG      �����  	 � � � �  Z@f9HH      �����   � � � �  n@g9II      �����   � � � �  i@h9JJ      �����  
 � � � �  n@i9KK      �����   � � � �    ~�n2
b`��$�� p"$�&�(              
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:� � �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@_ GG      �����   � � � �  d@` HH      �����   � � � �  d@` II      �����   � � � �  i@b JJ      �����   � � � �  Z@T <<      �����  � � � �  i@W'==      �����  � � � �  i@Y'>>      �����  � � � �  d@Z'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b���b!b&�,H3`4�6�7;    
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�P~ �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@f9GG      �����   � � � �  i@f9HH      �����   � � � �  _@h9II      �����   � � � �  n@h9JJ      �����   � � � �  L@Z9<<      �����  � � � �  d@[9==      �����  � � � �  i@\9>>      �����  � � � �  dA]9??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b���r��"�#�' ,�/    
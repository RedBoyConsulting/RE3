�?�?%�?5�?E�?T�?d�?u�?��?��?��?��?��?��?��?��?����������������!�����������������������������������������G��� �  �     ��   @  ����x��@�  ��������n��@�  �������� Z@N9<<      �����   � � � �  d@O9==      �����   � � � �  _@P9>>      �����   � � � �  _@Q9??      �����   � � � �  i@R9@@      �����   � � � �  s@aAA      �����  
 � � � �  n@`9BB      �����  	 � � � �  _@a9CC      �����   � � � �  i@\ DD      �����   � � � �  s@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@e9GG      �����   � � � �  Z@f9HH      �����   � � � �  n@g9II      �����   � � � �  i@h9JJ      �����   � � � �  n@i9KK      �����   � � � �   A@H <<      �����  � � � �  A@H <<      �����  � � � �  2@I ==      �����  � � � �    �
H	Vj8���.,� �#�(N,�/�02        
��#�4�D�T�d�q����������������������������������������������������������������������������������������������� �  p  P  	   �� 	 	 @  ����	n��@�  ��������  U@N9<<      �����   � � � �   n@P9==      �����   � � � �   Z@P9>>      �����   � � � �   U@Q9??      �����   � � � �   x@R9@@      �����   � � � �   d@S9AA      �����   � � � �   d@Q9BB      �����   � � � �   F@[ CC      �����   � � � �   K@V9DD      �����  	 � � � �    ����B(�            
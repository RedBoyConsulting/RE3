B` 5` ����ea U���������������������������������B�������������������������������������������������������������������������pr          ��   @  ����d��@�  ��������   @S;;;      �����   � � � �   i@H <<      �����   � � � �  i@H <<      �����   � � � �  d@I ==      �����   � � � �  i@J >>      �����   � � � �  x@K ??      �����   � � � �  n@L @@      �����   � � � �    ^*f�N  
��$���S�3�A�d�t�������������������������������������������������������������������������������� p  @     ��   @  ����d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@e9GG      �����   � � � �  d@f9HH      �����   � � � �  d@f9II      �����   � � � �  d@h9JJ      �����   � � � �    8�	.,b��j��6"            
��%�5�E�T�d�u�����������������5�E�U�e�q�������������������������%�������������G�@e �  @     ��   @  ����x��@�  ��������n��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  i@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  i@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �   Z@Rm<<      �����  � � � �  Z@Rm<<      �����  � � � �  i@[9==      �����  � � � �  x@\9>>      �����  � � � �  x@Y'??      ����� 	 � � � �  n@^'@@      ����� 
 � � � �  n@_9AA      �����  � � � �  2@N BB      �����  � � � �    8�TV
���z2\�P�| x$�%b'l*x+�,              
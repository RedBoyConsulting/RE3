��+�5�A�T�k�|���������������������������������������������������������������������������������@\ P  0     ��   @  ����d��@�  ��������  U@N9<<      �����   � � � �   P@K9==      �����   � � � �   @Cm>>      �����_   � � � �   @DF??      �����_   � � � �   F@R9@@      �����   � � � �   x@DFAA      �����_   � � � �   @MXBB      �����_   � � � �   @NZCC      �����_   � � � �   d@\9DD      �����   � � � �   <@X9EE      �����  	 � � � �   P@b FF      �����   � � � �   x@Y9GG      �����   � � � �   A@T HH      �����  
 � � � �   F@U II      �����   � � � �   P@X JJ      �����   � � � �   d@c KK      �����   � � � �   $@`��`�Z8 �!�"$n&�'�+
��$�>�D�T�c�t���������������t��������������������������������������������������������������������P P  0     ��   @  ����n��@�  �������� P@N9<<      �����   � � � �  Z@O9==      �����   � � � �  Z@P9>>      �����   � � � �  n@Um??      �����   � � � �  n@P9@@      �����   � � � �  Z@S9AA      �����   � � � �  Z@T9BB      �����  	 � � � �  @W9CC      �����   � � � �  n@V9DD      �����   � � � �  @W9EE      �����  
 � � � �  Z@^ FF      �����   � � � �  K@Y9GG      �����   � � � �  _@Z9HH      �����   � � � �   @S;II      �����   � � � �   @S;JJ      �����   � � � �  n@]9KK      �����   � � � �    ��������&%8(*  
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�p� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  _@f9GG      �����   � � � �  d@h9HH      �����   � � � �  Z@h9II      �����   � � � �  i@h9JJ      �����   � � � �  P@X'<<      �����  � � � �  d@W'==      �����  � � � �  d@X'>>      �����  � � � �  i@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,bJR�� $#J$�'r)->1N4    
 � %� 5� E� S�? c�? s�? ��? ��? ��?���� � ������ �g  ��P�    �     ��   @  ����d��@�  ��������  x@Qm;;      �����   � � � �   i@Rm<<      �����  	 � � � �   n@Sm==      �����   � � � �   n@Tm>>      �����  
 � � � �   n@Y'??      �����   � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �    @S;DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   A@T HH      �����M   � � � �    Z �<�x	V
�@l�      
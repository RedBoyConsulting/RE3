B` 5` ����ea U���������������������������������B��������������������������������������������������������������������������l          ��   @  ����d��@�  ��������   @S;;;      �����   � � � �   P@H <<      �����   � � � �  P@H <<      �����   � � � �  d@I ==      �����   � � � �  s@J >>      �����   � � � �  x@K ??      �����   � � � �  n@L @@      �����   � � � �    � 
�X�  
��������������������������������������*�������������������$���S�3�A�d�t���������������Pa �  P     ��   @  ����x��@�  ��������d��@�  ��������  �� �  ��������  i@Z9<<      �����   � � � �   x@[9==      �����   � � � �   Z@\9>>      �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  A@V'<<      ����� 	 � � � �  <@W'==      ����� 
 � � � �  @Tm>>      �����  � � � �  s@Q9??      �����  � � � �  Z@X @@      �����  � � � �  Z@]9KK      �����  � � � �  d@Y AA      �����  � � � �  @Z BB      �����  � � � �  d@[ CC      �����  � � � �  @\ DD      �����  � � � �  @[mEE      �����  � � � �  n@c FF      �����  � � � �  Z@e9GG      �����  � � � �  d@f9HH      �����  � � � �  d@g9II      �����  � � � �  U@h9JJ      �����  � � � �    8�	.,b��X"d$&"(*,      
��$���S�3�A�d�t���������������5�E�U�e�q�������������������������%�������������G�Pf �  P     ��   @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@Z9<<      �����   � � � �  7@Z9==      �����   � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@a9CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@f9GG      �����  	 � � � �  i@f9HH      �����  
 � � � �  _@h9II      �����   � � � �  n@h9JJ      �����   � � � �   Z@H <<      �����  � � � �  Z@H <<      �����  � � � �  d@[9==      �����  � � � �  s@\9>>      �����  � � � �  s@]9??      �����  � � � �  i@^9@@      �����  � � � �  i@_9AA      �����  � � � �  2@N BB      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    822���
 ������Z@>"n#�%�'�+�,
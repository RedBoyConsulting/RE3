B` 5` ����ea U���������������������������������B��������������������������������������������������������������������������n          ��   @  ����d��@�  ��������   @S;;;      �����   � � � �   x@H <<      �����   � � � �  x@H <<      �����   � � � �  d@I ==      �����   � � � �  i@H >>      �����   � � � �  x@K ??      �����   � � � �  n@L @@      �����   � � � �    ^��,�  
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�P� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  U@b GG      �����   � � � �  d@c HH      �����   � � � �  d@d II      �����   � � � �  i@d JJ      �����   � � � �  U@U'<<      �����  � � � �  _@W'==      �����  � � � �  _@X'>>      �����  � � � �  _@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b�F�� �"'�-�2�3J7    
��������������������������������������*�������������������$���S�3�A�d�t���������������� p  @     ��   @  ����x��@�  ��������s��@�  ��������  i@Z9<<      �����   � � � �   x@[9==      �����   � � � �   Z@\9>>      �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  K@V'<<      �����  � � � �  F@W'==      �����  � � � �  @Tm>>      �����  � � � �  _@U9??      �����  � � � �  _@X @@      �����  � � � �  _@S9AA      �����  � � � �    @S;BB      �����  � � � �    @S;CC      �����  � � � �  n@[ DD      �����  � � � �  @\ EE      �����  � � � �  @[mFF      ����� 	 � � � �  n@c GG      ����� 
 � � � �  Z@g9HH      �����  � � � �  Z@g9II      �����  � � � �  Z@i9JJ      �����  � � � �  x@i9KK      �����  � � � �    :lLt	 |��Z^��� �"            
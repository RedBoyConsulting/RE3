��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@f9GG      �����   � � � �  Z@f9HH      �����   � � � �  Z@h9II      �����   � � � �  x@h9JJ      �����   � � � �  U@U'<<      �����  � � � �  _@W'==      �����  � � � �  _@X'>>      �����  � � � �  _@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b�����#�$.(�)�,�/^4    
��������������������������������������*�������������������#�4�D�T�d�q���������������������������������  �  �  	   ��   @  ����x��@�  ��������	n��@�  ��������  i@Z9<<      �����  
 � � � �   x@[9==      �����   � � � �   Z@\9>>      �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   U@N9<<      �����  � � � �   n@P9==      �����  � � � �   Z@P9>>      �����  � � � �   U@Q9??      �����  � � � �   x@R9@@      �����  � � � �   d@S9AA      �����  � � � �   d@Q9BB      �����  � � � �   F@[ CC      �����  � � � �   K@V9DD      ����� 	 � � � �    ����B(����      
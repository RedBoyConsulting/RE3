B` %` 1�Ua ea Ea �������������������������������������������������������������������������������������������������������� x          ��   @  ����i��@�  ��������  s@C9<<      �����   � � � �  s@C9<<      �����   � � � �  d@I ==      �����   � � � �  F@J >>      �����   � � � �  Z@H ??      �����   � � � �  d@R9@@      �����   � � � �  (@M AA      �����   � � � �    � 	�� 
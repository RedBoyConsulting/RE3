��%�5�E�T�d�u���������������������������������������������������������������������������������� `  0     ��   @  ����x��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  i@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  i@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����  	 � � � �  Z@hHH      �����  
 � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �    8�TV
�h��0��z�!�"            
��%�5�E�T�d�u�������������������+�;�J�[�b�r��������������������������    �     ��   @  ����x��@�  ��������n��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  x@_AA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �   _@N9<<      �����  � � � �   n@T ==      ����� 	 � � � �   d@T>>      ����� 
 � � � �   n@W ??      �����  � � � �   n@\>@@      �����  � � � �   n@Y AA      �����  � � � �   i@\'BB      �����  � � � �   d@[ CC      �����  � � � �   P@V9DD      �����  � � � �   U@[mEE      �����  � � � �   i@^ FF      �����  � � � �   P@_ GG      �����  � � � �    8�TV

(�f� p!�"�#�$�(n+�/01�3\8�9b;=@A    
��%�5�E�T�d�u�������������������$���S�3�A�d�t����������������� �  @     ��    @  ����x��@�  ��������s��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  x@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �  K@V'<<      �����  � � � �  F@W'==      ����� 	 � � � �  @Tm>>      ����� 
 � � � �  _@U9??      �����  � � � �  _@X @@      �����  � � � �  _@S9AA      �����  � � � �    @S;BB      �����  � � � �    @S;CC      �����  � � � �  n@[ DD      �����  � � � �  @\ EE      �����  � � � �  @[mFF      �����  � � � �  n@c GG      �����  � � � �  i@i9HH      �����  � � � �  n@j9II      �����  � � � �  n@k9JJ      �����  � � � �  }@k9KK      �����  � � � �    8�TV
N�`�4���� �#�&�*R,�.~3�4�6&80;<<  
��%�5�E�����d�������������������������$���S�3�A�d�t���������������Ѓ �  @     ��    @  ����x��@�  ��������s��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �   @S;AA      �����   � � � �  s@`9BB      �����   � � � �   @S;CC      �����   � � � �   @S;DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �  K@V'<<      �����  � � � �  F@W'==      �����  � � � �  @Tm>>      �����  � � � �  _@U9??      ����� 	 � � � �  _@X @@      �����  � � � �  _@S9AA      ����� 	 � � � �    @S;BB      �����  � � � �    @S;CC      �����  � � � �  n@[ DD      ����� 
 � � � �  @\ EE      �����  � � � �  @[mFF      �����  � � � �  n@c GG      �����  � � � �  i@i9HH      �����  � � � �  n@h9II      �����  � � � �  s@j9JJ      �����  � � � �  n@k9KK      �����  � � � �    � �JH~�	��d����.�  #�')�*d,n/z0            
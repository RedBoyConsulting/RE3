��$���S�3�A�d�t�������������������������������!�����������������������������������������G�`T �  P     ��   @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  U@c'GG      �����   � � � �  Z@d'HH      �����   � � � �  d@d'II      �����   � � � �  _@d'JJ      �����   � � � �   Z@H <<      �����  � � � �  Z@H <<      �����  � � � �  2@I ==      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,bVH�!>#d$�'\)�*        
��*�2�A�Q�j�����������������������������������������������������'"�����������������������������������������g���  �  �     �� 
 
 @  ����d��@�  ��������d��@�  ��������  d@I<<      �����   � � � �   d@M>==      �����   � � � �   d@K>>      �����   � � � �   d@O>??      �����   � � � �   d@R9@@      �����   � � � �   d@S9AA      �����   � � � �   d@Q6BB      �����   � � � �   -
H <<      ����� 	 � � � �   -
H <<      ����� 	 � � � �   
I ==      ����� 
 � � � �    �t*�4����          
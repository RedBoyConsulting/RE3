��������������������������������������*�������������������"�;�D�S�b�s���������������t���{ p  @     ��   @  ����x��@�  ��������n��@�  ��������  i@Z9<<      �����   � � � �   x@[9==      �����   � � � �   Z@^>>      �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  P@T <<      ����� 
 � � � �  Z@U ==      �����  � � � �  Z@P9>>      �����  � � � �  n@Um??      �����  � � � �  n@P9@@      �����  � � � �  Z@S9AA      �����  � � � �  Z@T9BB      �����  � � � �  x@W9CC      �����  � � � �  n@V9DD      �����  � � � �  @W9EE      �����  � � � �  n@d9FF      �����  � � � �  K@Y9GG      ����� 	 � � � �  _@Z9HH      �����  � � � �    @S;II      �����  � � � �    @S;JJ      �����  � � � �  n@]9KK      �����  � � � �    :z(�	nL�D$�#�%�'�)�+b/            
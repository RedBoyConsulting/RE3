��%�5�E�T�d�u�������������������*�2�A�Q�j�������������������������������������@� `        ��   @  ����x��@�  ��������n��@�  �������� d@Z9<<      �����   � � � �  i@[9==      �����   � � � �  _@\9>>      �����   � � � �  i@]9??      �����   � � � �  x@^9@@      �����   � � � �  i@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  i@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@gGG      �����  	 � � � �  Z@hHH      �����  
 � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �  d@I<<      �����  � � � �  d@M>==      �����  � � � �  d@K>>      �����  � � � �  d@O>??      �����  � � � �  d@R9@@      �����  � � � �  d@S9AA      �����  � � � �  d@Q6BB      �����  � � � �    8�TV
�h��0��z�!�"J'�)�.r1�25(:              
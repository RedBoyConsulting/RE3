��$���S�3�A�d�t�������������������������������������������������������������������������������U p  @     ��   @  ����d��@�  ��������  �� �  �������� F@N9<<      �����   � � � �  <@W'==      �����  	 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����  
 � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@` GG      �����   � � � �  d@a HH      �����   � � � �  d@b II      �����   � � � �  n@d JJ      �����   � � � �    8�	.d��.�\$�%�(�*            
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  U@` GG      �����   � � � �  n@a HH      �����   � � � �  i@a II      �����   � � � �  i@b JJ      �����   � � � �  d@U <<      �����  � � � �  d@V ==      �����  � � � �  d@W >>      �����  � � � �  i@Y ??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b�����$�%&+�2T9z:�=    
��$���S�3�A�d�t���������������5�E�U�e�q�������������������������%�������������G���  �  P     ��   @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@V'<<      �����   � � � �  <@W'==      �����   � � � �   @S;>>      �����   � � � �   @S;??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �   @S;AA      �����   � � � �   @S;BB      �����   � � � �   @S;CC      �����   � � � �   @S;DD      �����   � � � �   @S;EE      �����   � � � �   @S;FF      �����   � � � �  d@f9GG      �����   � � � �  i@f9HH      �����   � � � �  _@h9II      �����   � � � �  n@h9JJ      �����  	 � � � �   Z@H <<      ����� 
 � � � �  Z@H <<      ����� 
 � � � �  d@[9==      �����  � � � �  s@\9>>      �����  � � � �  s@]9??      �����  � � � �  i@^9@@      �����  � � � �  i@_9AA      �����  � � � �  2@N BB      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    ��B	����|b6`�              
��������������������������������������*�������������������"�3�B�R�b�r���������������������������`�           ��   @  ����x��@�  ��������i��@�  ��������  i@Z9<<      �����   � � � �   x@[9==      �����   � � � �   Z@\9>>      �����   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  2@N9<<      �����  � � � �  @O9==      �����  � � � �  Z@P9>>      �����  � � � �  @Um??      �����  � � � �  @R9@@      �����  � � � �  s@S9AA      �����  � � � �  @T9BB      �����  � � � �  n@U9CC      ����� 	 � � � �  <@V9DD      �����  � � � �  F@W9EE      �����  � � � �  (@X9FF      ����� 
 � � � �    � �v0���r����    
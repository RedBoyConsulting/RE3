��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@a'GG      �����   � � � �  d@c'HH      �����   � � � �  d@b'II      �����   � � � �  d@d'JJ      �����   � � � �  Z@V'<<      �����  � � � �  Z@U ==      �����  � � � �  d@X'>>      �����  � � � �  Z@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b�~�*�$l&|+20�6�7;    
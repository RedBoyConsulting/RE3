��%�5�E�T�d�u���������������������������������������������������������������������������������`< `  0     ��   @  ����x��@�  �������� _@T <<      �����   � � � �  i@O9==      �����   � � � �  d@V >>      �����  
 � � � �  n@W ??      �����  	 � � � �  n@R9@@      �����   � � � �  x@aAA      �����   � � � �  s@`9BB      �����   � � � �  i@f;CC      �����   � � � �  n@b9DD      �����   � � � �  x@f EE      �����   � � � �  x@i;FF      �����   � � � �  d@g9GG      �����   � � � �  Z@hHH      �����   � � � �  n@iII      �����   � � � �  i@jJJ      �����   � � � �  n@kKK      �����   � � � �    ~��
�
�T�����` �"�'            
��-�=�N�_�c���}�����������������������������������������������������������������������������������������p\ �  �     ��   @  ����x��@�  ��������  Z@Rm<<      �����   � � � �   d@V9==      �����   � � � �   n@\9>>      �����   � � � �   s@W ??      �����   � � � �   s@R9@@      �����   � � � �   x@['AA      �����  
 � � � �   n@e;BB      �����   � � � �   n@[9CC      �����   � � � �   d@_9DD      �����O   � � � �   n@d9FF      �����   � � � �   d@j GG      �����  	 � � � �    *��f( X#)�+        
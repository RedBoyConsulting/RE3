�?�?+�?;�?J�?[�?b�?r�?��?��?��?��?��������������������������������'"�����������������������������������������g�� @        ��   @  ����d��@�  ��������n��@�  ��������  _@N9<<      �����   � � � �   n@T ==      �����   � � � �   d@T>>      �����   � � � �   n@U;??      �����   � � � �   n@\>@@      �����   � � � �   n@Y AA      �����   � � � �   i@\'BB      �����   � � � �   d@[ CC      �����   � � � �   P@V9DD      �����   � � � �   U@\mFF      �����  	 � � � �   i@_ GG      �����  
 � � � �   P@_;HH      �����N   � � � �   -
H <<      �����  � � � �   -
H <<      �����  � � � �   
I ==      �����  � � � �    �x	j�.FT��B r!
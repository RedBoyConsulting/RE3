��+�5�A�T�k�|����������������������������������������������������������������������������������� M 0       ��   @  ����d��@�  �������� d@EF<<      �����_   � � � �  P@A ==      �����_   � � � �  @Cm>>      �����_   � � � �  @DF??      �����_   � � � �  A@L @@      �����   � � � �  x@DFAA      �����_   � � � �  @MXBB      �����_   � � � �  @NZCC      �����_   � � � �  d@\9DD      �����   � � � �  <@X9EE      �����   � � � �  P@b FF      �����  	 � � � �  }@[9GG      �����   � � � �  A@T HH      �����   � � � �  F@U II      �����  
 � � � �  P@X JJ      �����   � � � �   2V
r�0�
 h"6#�$0&'v(�)  
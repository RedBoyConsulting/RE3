��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:�p� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@b'GG      �����   � � � �  d@b'HH      �����   � � � �  d@c'II      �����   � � � �  Z@e'JJ      �����   � � � �  U@W'<<      �����  � � � �  Z@X'==      �����  � � � �  d@Y'>>      �����  � � � �  d@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b���B�#�$L*�0�6�7.;    
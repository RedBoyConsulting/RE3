��$���S�3�A�d�t������������������������������������������������������������������������������� I p  @     ��   @  ����d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@a'GG      �����   � � � �  d@c'HH      �����   � � � �  d@b'II      �����   � � � �  d@d'JJ      �����   � � � �    8�	.,b�~�*�$�%$)            
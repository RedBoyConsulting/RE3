��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:� w �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  Z@f9GG      �����   � � � �  Z@f9HH      �����   � � � �  Z@h9II      �����   � � � �  x@h9JJ      �����   � � � �  _@[9<<      �����  � � � �  d@^9==      �����  � � � �  Z@\9>>      �����  � � � �  i@^9??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b��j��6"$�'�+�.    
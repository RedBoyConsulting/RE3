��$���S�3�A�d�t�������������������������������!�����������������������������������������G�`9 �  P     ��   @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@e9GG      �����   � � � �  d@f9HH      �����   � � � �  d@g9II      �����   � � � �  d@g9JJ      �����   � � � �   s@N9<<      �����  � � � �  s@N9<<      �����  � � � �  <@I ==      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b��Z���#L$,'        
��$���S�3�A�d�t�����������������$���S�3�A�d�t���������+�:��� �  P     ��   @  ����d��@�  ��������d��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  U@c'GG      �����   � � � �  Z@d'HH      �����   � � � �  d@d'II      �����   � � � �  _@d'JJ      �����   � � � �  P@X'<<      �����  � � � �  d@W'==      �����  � � � �  d@X'>>      �����  � � � �  i@Y'??      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,bVH�!�!'�,�2�4�5T9    
��$�>�D�T�c���������������t��������������������������������������������������������������������R `  0     ��   @  ����n��@�  �������� P@T <<      �����  
 � � � �  Z@U ==      �����   � � � �  Z@P9>>      �����   � � � �  n@Um??      �����   � � � �  n@P9@@      �����   � � � �  Z@S9AA      �����   � � � �  Z@T9BB      �����   � � � �  x@W9CC      �����   � � � �  n@V9DD      �����   � � � �  @W9EE      �����   � � � �  n@d9FF      �����   � � � �  K@Y9GG      �����  	 � � � �  _@Z9HH      �����   � � � �  Z@a II      �����   � � � �  d@b JJ      �����   � � � �  n@]9KK      �����   � � � �    :z(�	nL�D$�#�%�'x(R*              
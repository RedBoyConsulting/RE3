 � %� 5� E� S�? c�? s�? ��? ��? ��?���� � ������ �g  ��`�    �     ��   @  ����d��@�  ��������  x@Qm;;      �����   � � � �   s@T <<      �����  
 � � � �   n@U ==      �����   � � � �   n@V >>      �����   � � � �   x@Y'??      �����  	 � � � �  7@L @@      �����   � � � �  U@M AA      �����   � � � �  Z@T9BB      �����   � � � �  K@[ CC      �����   � � � �    @S;DD      �����   � � � �    @S;::      �����   � � � �    @S;::      �����   � � � �  d@\9GG      �����_   � � � �   A@T HH      �����M   � � � �    Z �<�x	

����      
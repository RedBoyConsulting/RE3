��$���S�3�A�d�t���������������5�E�U�e�q�������������������������%�������������G��g �  P     �� !  @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  d@e9GG      �����   � � � �  d@f9HH      �����   � � � �  d@g9II      �����   � � � �  d@g9JJ      �����   � � � �   Z@Rm<<      �����  � � � �  Z@Rm<<      �����  � � � �  d@[9==      �����  � � � �  s@\9>>      �����  � � � �  s@]9??      �����  � � � �  i@^9@@      �����  � � � �  i@_9AA      �����  � � � �  2@N BB      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b��Z���#�#�$j%>&h)�+�,              
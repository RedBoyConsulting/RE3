��*�2�A�Q�j������������������������������������������������������������������������������������������������������  0       ��   @  ����d��@�  ��������  d@I<<      �����   � � � �   d@M>==      �����   � � � �   d@K>>      �����   � � � �   d@O>??      �����   � � � �   d@R9@@      �����   � � � �   d@S9AA      �����   � � � �   d@Q6BB      �����   � � � �    �t*�4��              
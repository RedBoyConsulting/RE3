��$���S�3�A�d�t�������������������������������!�����������������������������������������G� [ �  P     ��   @  ����d��@�  ��������n��@�  ��������  �� �  �������� A@V'<<      �����  	 � � � �  <@W'==      �����  
 � � � �  @Tm>>      �����   � � � �  s@Q9??      �����   � � � �  Z@X @@      �����   � � � �  Z@]9KK      �����   � � � �  d@Y AA      �����   � � � �  @Z BB      �����   � � � �  d@[ CC      �����   � � � �  @\ DD      �����   � � � �  @[mEE      �����   � � � �  n@c FF      �����   � � � �  U@b'GG      �����   � � � �  _@b'HH      �����   � � � �  d@c'II      �����   � � � �  d@d'JJ      �����   � � � �   F@H <<      �����  � � � �  F@H <<      �����  � � � �  <@I ==      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    8�	.,b��6n�^$@*d+        